.title Parallel Resistors 
V1 N001 0 5
R1 N001 0 2
R2 N001 0 3

.control 
.option savecurrents 
dc V1 0 5 0.1 
plot @R1[i], @R2[i]
.endc

.end